`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:38:14 05/01/2025 
// Design Name: 
// Module Name:    mux_16b_8to1 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mux_16b_8to1(
    input [2:0]sel,
	 input [15:0]data0,data1,data2,data3,data4,data5,data6,data7,
	 output [15:0]out
    );
	
endmodule
